`timescale 1ns / 1ps
module t_test;
  reg clk,rst,start;
  reg [0:323]sudoku_given;
  wire completed;
  wire [0:323] sudoku_out;
 candidate_type1     m1(completed,sudoku_out,rst,start,clk,sudoku_given);
  initial
    begin
     rst=1'b0;
      start=1'b0;
       #8 rst=1'b1;
      #152 rst=1'b0;
      #1 sudoku_given=324'h735468912064139058819527463978613524126954837453782196342891675681275349097346081;//001957063000806070769130805007261350312495786056378000108609507090710608674583000;//286045700709130506031006400908000204120600075000400601850200000000709300000080000;
      #1 start=1'b1;
      #10 @(completed)
      $display($time);
       #5 $write("%81h",sudoku_out);
      #10 $finish;
      end  
  initial
    begin
      clk=1'b0;
      forever
        #5 clk=~clk;
    end
endmodule
  //546971203972836510801452967000305600765140308029768451053684702094217835280590146
  //546971283972836514831452967418325679765149328329768451153684792694217835287593146
//281957463435826971769134825847261359312495786956378214128649537593712648674583192